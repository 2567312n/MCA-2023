BZh91AY&SY�� J_�Ryg������?���    ��  �    =M�OP � ��� =C@4EOP�2 hh4 P    8ɓF!��hbh�& da4i�d�2h�4��MMd��&�4���&M��	���L����Ѧ�A�I� &� L&��<P44d���6�P�*P�̓C����`$�I$��'�~o��L!��md���c���.��U'�M?�C�K4��5nf���iۂ���I¶P���KT��d�I�!qI����V��F�q�bT5T��;m�n���|�m��[Vzz���k�V���Svkc=1����獻%Mp�ޛ|�b�ae�Z�챞���-e�ulƯjzK~yɁ�a��u^��SJ��/c���Ɍ�k�]�\�N�ɔo�Z޷t�#,zL�`�8�$��F3\N�g:�Rv4{W7ft^�~�F�ιq���ڢ����D�r�a��iƛ(�We��}�-J��?S��,Tʾvl��LBֲ6�;��ZZ�K��:�MT�I���]05Ҟs<��ٔ�X��p�ݸ�����UQ�L�2l��d��ٙ��4b����:^c�������,�U�UUUUUU�eԴh����鞵M�~e�e�����Qn8F�K����Z�srYmn��)/'M�K�m5l,aQz��,ɹhgRh��UY�lڸ�+2�!�i����9)UUwiaTl\8�T!d�	L�$?#��m[����;#�)'Su�0U��Jj�P]D���k&�)�X��y5\�Ϲj��û���c��)���Oœ���y����6M���G8��A�)U0��s��bO���2�
��,�d\}Qˣ�o��7�Ruln������u���'��b��N3sΧll#k���W��g��e�u�N�)^i͠�h�ix�W��T�dT�1�&;�"72�z%�K_@�Lϻ��(�1b������G�4�t��Q����yIx����z)����J���/�]��l�0���i%����M�̩b��׃k"���N��>��v��B�X�$vm+'!�̋��G��!d{-[�e7�>��wI�6O���:~9;�dN���KvCr�%�q��Z=��<�ں�)R��z�����R���b�˽���(Е��1�o��|�[��.�ɱ�5Y֔�b�c'�O�Yuۤ�G)�W�q�3��:�iį1�*}����h�]�'lģ�B���4%��g�Ѻ|d��	�y
Z�9c5h�����5��38��,?���9�����(��)R�)��	�R<�ĩ��3�4���^bco��ub�s8��Z�V��yV,Y;%%��"nݤh��k�%-E�H��?0��TѤ���F�&���i!^G�V�R_��=��FsT<���d÷�'7�7C{�6�{���s.G�'V����:�w�eXy��'���骴���%�k�{�5�g'��N�(�p��w���QH��C�=�����F�����R��6����Ŝ��¡Vw�Z�<�cee%�a]/5��Y��wywbŨ�^I�����U}ծ�N�G3��G7	����<���5j�&�rTp�m��<��h�Ͱfa�XE�94H����>�Qdtz��K�Q�Q�zv6���]��sՄ���u���RM���.�:;�g�S���8�)�
UA�L
Rc�LF��_��|��.�p�!
-8