BZh91AY&SY~e� HߩRyg������?���    ��  �    �4���4   ��  �MC�F�  ��   �&M��	���L����Ѧ�A�dɣ�C414i�20�4�2c��4bh`&�&�2bFF�aL$@@�Bdhi�FBOQ�����:�JyRh5Ќ�I$�XD����[�c�d��k����U~O�7�?��_KFo3���>�;�]6?R�p��-*A�KP�l�%�Li�MWXd��j��TmWF%CUH��چ����p���`�j�OTx�{�F��_�Mذi��4Ɨ�%���l��U�Ϟ,[l,���E6u��[//ڵ�YҰ������3����Y����L*�tv=n��Lf}�����﬙G
��l}�1á��#�RH9��k���l�U��#ع�3��zz��
���s�t�&�nQIJ���b3�a���q�T��vg��,r��2����%�����UF

�kZCZ�EH]�Z�Գ�UcI��G���5�j:���u]�/|�˖�v����g�*����f80��yK⶧��F��6z<�ӭc��'j��,�U�UUUUUU�
��Z4z<G��y�SmߙtYz�{>��Qn8F�K��6]��ZT{jכi,�/���SR��v�f�]/Q\�nZԙ��UVh�6�6J̣EHaZm���9)UUwiaTlذ��PZR�'���z���.�q��pDdf�CI�M�kk@\�"@s< btG#����s$�`)�X��x�\�Ϲj��û���c��źL;7�6�N�c����Q��c�)J�n��P��'��2�
��2�,��lr��8?��|�{c�dG�|郺����e�iw'�槊6���I�ګ����˩u�?��,��x>MK�R�-�M����1�&<"72�z%�|�af}�v,7bQbŃc;qh������{NP�����K����=3��t����*����+:�H���_-$����)�ٕ,^^z�mdSV3i�Gϔa���cV��w�nҷ�r��̻��f|d�#���p���f��R�)�&,�=��Q���a�z��u��-����;�Z=��;ѵu*R�<���y�R���b������(МS'��רz�,�m��1��ħsŌ�Gd��e�n��9O*�;����6��#N%yN��ߛ=F����|!I☔tP���Ƅ��)���T��]���;�Z�9e5~�]�H��`��|s0#��a���d2N�,�j��)��T��l�`T�	bT�o)њIRR/11��杘���������oZT^��bŪ�S�R[H���+q��IE�F�R-f��(hi�j�F;%�*��09<��פ�x��[L]�����3���P�JPo��f؟���.m��m|JN�������M�n�E�P{���E�a�$�\=5V����w���ػ���r�%Rtb��%Ț�E"����O���j���2�08	��le�,�g(�
���k�����Z��府+7��&�X�k�4�����c}�����ٳ��#��ub(��2Ѵ��bqG�7��\��NJ���ۥ�yu�у�`��8���rh��{�P�������)0K��#�OFͭÁ�uE�YG=XL\�gY�ٙ�$�z�a�������utS���`R��:��n?���?�]��BA���D